`resetall
`timescale 1ns/1ns

module moore_fsm1_tb;
    reg Clock, Resetn, w;
    wire z;